module OR(
    input wire S1,
    input wire S2,
    output wire F
);

assign F = S1|S2;

endmodule